../node/pkg.vhd