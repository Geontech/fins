--==============================================================================
-- Company:     Geon Technologies, LLC
-- Author:      Josh Schindehette
-- Copyright:   (c) 2019 Geon Technologies, LLC. All rights reserved.
--              Dissemination of this information or reproduction of this
--              material is strictly prohibited unless prior written
--              permission is obtained from Geon Technologies, LLC
-- Description: This is the top level testbench of the FINS test module
-- Reset Type:  Synchronous
--==============================================================================

-- Standard Libraries
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use ieee.math_real.all;
library std;
use std.textio.all;

-- User Libraries
library work;
use work.test_top_pkg.all;
use work.test_top_axilite_verify.all;
use work.test_middle_axilite_verify.all;
use work.test_bottom_swconfig_verify.all;

-- Entity
entity test_top_tb is
end entity test_top_tb;

-- Architecture
architecture rtl of test_top_tb is

  -- Device Under Test interface
  signal s_axis_myinput_tvalid  : std_logic;
  signal s_axis_myinput_tlast   : std_logic;
  signal s_axis_myinput_tdata   : std_logic_vector(PORTS_WIDTH-1 downto 0);
  signal m_axis_myoutput_tvalid : std_logic;
  signal m_axis_myoutput_tlast  : std_logic;
  signal m_axis_myoutput_tdata  : std_logic_vector(PORTS_WIDTH-1 downto 0);
  signal S_AXI_ACLK             : std_logic;
  signal S_AXI_ARESETN          : std_logic;
  signal S_AXI_AWADDR           : std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
  signal S_AXI_AWPROT           : std_logic_vector(2 downto 0);
  signal S_AXI_AWVALID          : std_logic;
  signal S_AXI_AWREADY          : std_logic;
  signal S_AXI_WDATA            : std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
  signal S_AXI_WSTRB            : std_logic_vector((PROPS_DATA_WIDTH/8)-1 downto 0);
  signal S_AXI_WVALID           : std_logic;
  signal S_AXI_WREADY           : std_logic;
  signal S_AXI_BRESP            : std_logic_vector(1 downto 0);
  signal S_AXI_BVALID           : std_logic;
  signal S_AXI_BREADY           : std_logic;
  signal S_AXI_ARADDR           : std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
  signal S_AXI_ARPROT           : std_logic_vector(2 downto 0);
  signal S_AXI_ARVALID          : std_logic;
  signal S_AXI_ARREADY          : std_logic;
  signal S_AXI_RDATA            : std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
  signal S_AXI_RRESP            : std_logic_vector(1 downto 0);
  signal S_AXI_RVALID           : std_logic;
  signal S_AXI_RREADY           : std_logic;
  signal S_AXI_MIDDLE_ACLK      : std_logic;
  signal S_AXI_MIDDLE_ARESETN   : std_logic;
  signal S_AXI_MIDDLE_AWADDR    : std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
  signal S_AXI_MIDDLE_AWPROT    : std_logic_vector(2 downto 0);
  signal S_AXI_MIDDLE_AWVALID   : std_logic;
  signal S_AXI_MIDDLE_AWREADY   : std_logic;
  signal S_AXI_MIDDLE_WDATA     : std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
  signal S_AXI_MIDDLE_WSTRB     : std_logic_vector((PROPS_DATA_WIDTH/8)-1 downto 0);
  signal S_AXI_MIDDLE_WVALID    : std_logic;
  signal S_AXI_MIDDLE_WREADY    : std_logic;
  signal S_AXI_MIDDLE_BRESP     : std_logic_vector(1 downto 0);
  signal S_AXI_MIDDLE_BVALID    : std_logic;
  signal S_AXI_MIDDLE_BREADY    : std_logic;
  signal S_AXI_MIDDLE_ARADDR    : std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
  signal S_AXI_MIDDLE_ARPROT    : std_logic_vector(2 downto 0);
  signal S_AXI_MIDDLE_ARVALID   : std_logic;
  signal S_AXI_MIDDLE_ARREADY   : std_logic;
  signal S_AXI_MIDDLE_RDATA     : std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
  signal S_AXI_MIDDLE_RRESP     : std_logic_vector(1 downto 0);
  signal S_AXI_MIDDLE_RVALID    : std_logic;
  signal S_AXI_MIDDLE_RREADY    : std_logic;
  signal s_swconfig_clk         : std_logic;
  signal s_swconfig_reset       : std_logic;
  signal s_swconfig_address     : std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
  signal s_swconfig_wr_enable   : std_logic;
  signal s_swconfig_wr_data     : std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
  signal s_swconfig_rd_enable   : std_logic;
  signal s_swconfig_rd_valid    : std_logic;
  signal s_swconfig_rd_data     : std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);

  -- Testbench
  signal simulation_done  : boolean := false;
  constant AXI_CLK_PERIOD : time := 5 ns;
  signal myinput_enable   : std_logic := '0';

begin

  -- Connect the AXI clocks and resets
  S_AXI_MIDDLE_ACLK    <= S_AXI_ACLK;
  S_AXI_MIDDLE_ARESETN <= S_AXI_ARESETN;

  -- Device Under Test
  u_dut : entity work.test_top
    port map (
      s_axis_myinput_tvalid  => s_axis_myinput_tvalid  ,
      s_axis_myinput_tlast   => s_axis_myinput_tlast   ,
      s_axis_myinput_tdata   => s_axis_myinput_tdata   ,
      m_axis_myoutput_tvalid => m_axis_myoutput_tvalid ,
      m_axis_myoutput_tlast  => m_axis_myoutput_tlast  ,
      m_axis_myoutput_tdata  => m_axis_myoutput_tdata  ,
      S_AXI_ACLK             => S_AXI_ACLK             ,
      S_AXI_ARESETN          => S_AXI_ARESETN          ,
      S_AXI_AWADDR           => S_AXI_AWADDR           ,
      S_AXI_AWPROT           => S_AXI_AWPROT           ,
      S_AXI_AWVALID          => S_AXI_AWVALID          ,
      S_AXI_AWREADY          => S_AXI_AWREADY          ,
      S_AXI_WDATA            => S_AXI_WDATA            ,
      S_AXI_WSTRB            => S_AXI_WSTRB            ,
      S_AXI_WVALID           => S_AXI_WVALID           ,
      S_AXI_WREADY           => S_AXI_WREADY           ,
      S_AXI_BRESP            => S_AXI_BRESP            ,
      S_AXI_BVALID           => S_AXI_BVALID           ,
      S_AXI_BREADY           => S_AXI_BREADY           ,
      S_AXI_ARADDR           => S_AXI_ARADDR           ,
      S_AXI_ARPROT           => S_AXI_ARPROT           ,
      S_AXI_ARVALID          => S_AXI_ARVALID          ,
      S_AXI_ARREADY          => S_AXI_ARREADY          ,
      S_AXI_RDATA            => S_AXI_RDATA            ,
      S_AXI_RRESP            => S_AXI_RRESP            ,
      S_AXI_RVALID           => S_AXI_RVALID           ,
      S_AXI_RREADY           => S_AXI_RREADY           ,
      S_AXI_MIDDLE_ACLK      => S_AXI_MIDDLE_ACLK      ,
      S_AXI_MIDDLE_ARESETN   => S_AXI_MIDDLE_ARESETN   ,
      S_AXI_MIDDLE_AWADDR    => S_AXI_MIDDLE_AWADDR    ,
      S_AXI_MIDDLE_AWPROT    => S_AXI_MIDDLE_AWPROT    ,
      S_AXI_MIDDLE_AWVALID   => S_AXI_MIDDLE_AWVALID   ,
      S_AXI_MIDDLE_AWREADY   => S_AXI_MIDDLE_AWREADY   ,
      S_AXI_MIDDLE_WDATA     => S_AXI_MIDDLE_WDATA     ,
      S_AXI_MIDDLE_WSTRB     => S_AXI_MIDDLE_WSTRB     ,
      S_AXI_MIDDLE_WVALID    => S_AXI_MIDDLE_WVALID    ,
      S_AXI_MIDDLE_WREADY    => S_AXI_MIDDLE_WREADY    ,
      S_AXI_MIDDLE_BRESP     => S_AXI_MIDDLE_BRESP     ,
      S_AXI_MIDDLE_BVALID    => S_AXI_MIDDLE_BVALID    ,
      S_AXI_MIDDLE_BREADY    => S_AXI_MIDDLE_BREADY    ,
      S_AXI_MIDDLE_ARADDR    => S_AXI_MIDDLE_ARADDR    ,
      S_AXI_MIDDLE_ARPROT    => S_AXI_MIDDLE_ARPROT    ,
      S_AXI_MIDDLE_ARVALID   => S_AXI_MIDDLE_ARVALID   ,
      S_AXI_MIDDLE_ARREADY   => S_AXI_MIDDLE_ARREADY   ,
      S_AXI_MIDDLE_RDATA     => S_AXI_MIDDLE_RDATA     ,
      S_AXI_MIDDLE_RRESP     => S_AXI_MIDDLE_RRESP     ,
      S_AXI_MIDDLE_RVALID    => S_AXI_MIDDLE_RVALID    ,
      S_AXI_MIDDLE_RREADY    => S_AXI_MIDDLE_RREADY    ,
      s_swconfig_clk         => s_swconfig_clk         ,
      s_swconfig_reset       => s_swconfig_reset       ,
      s_swconfig_address     => s_swconfig_address     ,
      s_swconfig_wr_enable   => s_swconfig_wr_enable   ,
      s_swconfig_wr_data     => s_swconfig_wr_data     ,
      s_swconfig_rd_enable   => s_swconfig_rd_enable   ,
      s_swconfig_rd_valid    => s_swconfig_rd_valid    ,
      s_swconfig_rd_data     => s_swconfig_rd_data     
    );

  -- File input/output streams
  -- NOTE: The source/sink filepaths are relative to where the simulation is executed
  u_file_io : entity work.test_top_streams
    generic map (
      G_MYINPUT_SOURCE_FILEPATH => "../../../../../../sim_data/sim_source_myinput.txt",
      G_MYOUTPUT_SINK_FILEPATH  => "../../../../../../sim_data/sim_sink_myoutput.txt"
    )
    port map (
      simulation_done        => simulation_done,
      m_axis_myinput_clk     => S_AXI_ACLK,
      m_axis_myinput_enable  => myinput_enable,
      m_axis_myinput_tdata   => s_axis_myinput_tdata,
      m_axis_myinput_tvalid  => s_axis_myinput_tvalid,
      m_axis_myinput_tlast   => s_axis_myinput_tlast,
      m_axis_myinput_tready  => '1',
      s_axis_myoutput_clk    => S_AXI_ACLK,
      s_axis_myoutput_tdata  => m_axis_myoutput_tdata,
      s_axis_myoutput_tvalid => m_axis_myoutput_tvalid,
      s_axis_myoutput_tlast  => m_axis_myoutput_tlast,
      s_axis_myoutput_tready => open
    );

  -- AXI Clock
  w_axi_clk : process
  begin
    if (simulation_done = false) then
      S_AXI_ACLK <= '0';
      s_swconfig_clk <= '0';
      wait for AXI_CLK_PERIOD/2;
      S_AXI_ACLK <= '1';
      s_swconfig_clk <= '1';
      wait for AXI_CLK_PERIOD/2;
    else
      wait;
    end if;
  end process w_axi_clk;


  w_test_procedure : process
    variable my_line : line;
  begin

    --**************************************************
    -- Reset
    --**************************************************
    S_AXI_ARESETN <= '0';
    s_swconfig_reset <= '1';
    wait for AXI_CLK_PERIOD*10;
    S_AXI_ARESETN <= '1';
    s_swconfig_reset <= '0';
    if (S_AXI_ARESETN = '0') then
      wait until (S_AXI_ARESETN = '1');
    end if;

    --**************************************************
    -- Verify registers
    --**************************************************
    test_top_axilite_verify (
      S_AXI_ACLK,
      S_AXI_ARESETN,
      S_AXI_AWADDR,
      S_AXI_AWPROT,
      S_AXI_AWVALID,
      S_AXI_AWREADY,
      S_AXI_WDATA,
      S_AXI_WSTRB,
      S_AXI_WVALID,
      S_AXI_WREADY,
      S_AXI_BRESP,
      S_AXI_BVALID,
      S_AXI_BREADY,
      S_AXI_ARADDR,
      S_AXI_ARPROT,
      S_AXI_ARVALID,
      S_AXI_ARREADY,
      S_AXI_RDATA,
      S_AXI_RRESP,
      S_AXI_RVALID,
      S_AXI_RREADY
    );

    --**************************************************
    -- Verify registers for test_middle module
    --**************************************************
    test_middle_axilite_verify (
      S_AXI_MIDDLE_ACLK,
      S_AXI_MIDDLE_ARESETN,
      S_AXI_MIDDLE_AWADDR,
      S_AXI_MIDDLE_AWPROT,
      S_AXI_MIDDLE_AWVALID,
      S_AXI_MIDDLE_AWREADY,
      S_AXI_MIDDLE_WDATA,
      S_AXI_MIDDLE_WSTRB,
      S_AXI_MIDDLE_WVALID,
      S_AXI_MIDDLE_WREADY,
      S_AXI_MIDDLE_BRESP,
      S_AXI_MIDDLE_BVALID,
      S_AXI_MIDDLE_BREADY,
      S_AXI_MIDDLE_ARADDR,
      S_AXI_MIDDLE_ARPROT,
      S_AXI_MIDDLE_ARVALID,
      S_AXI_MIDDLE_ARREADY,
      S_AXI_MIDDLE_RDATA,
      S_AXI_MIDDLE_RRESP,
      S_AXI_MIDDLE_RVALID,
      S_AXI_MIDDLE_RREADY
    );

    --**************************************************
    -- Verify registers for test_bottom module
    --**************************************************
    test_bottom_swconfig_verify (
      s_swconfig_clk       ,
      s_swconfig_reset     ,
      s_swconfig_address   ,
      s_swconfig_wr_enable ,
      s_swconfig_wr_data   ,
      s_swconfig_rd_enable ,
      s_swconfig_rd_valid  ,
      s_swconfig_rd_data   
    );

    --**************************************************
    -- Process data
    --**************************************************
    myinput_enable <= '1';
    wait until falling_edge(m_axis_myoutput_tlast);

    --**************************************************
    -- End Simulation
    --**************************************************
    write(my_line, string'("***** SIMULATION PASSED *****"));
    writeline(output, my_line);
    simulation_done <= true;
    wait;

  end process w_test_procedure;

end rtl;
