--==============================================================================
-- Company:     Geon Technologies, LLC
-- Author:      Josh Schindehette
-- Copyright:   (c) 2019 Geon Technologies, LLC. All rights reserved.
--              Dissemination of this information or reproduction of this
--              material is strictly prohibited unless prior written
--              permission is obtained from Geon Technologies, LLC
-- Description: This is the top level of the FINS test module
-- Reset Type:  Synchronous
--==============================================================================

-- Standard Libraries
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

-- User Libraries
library work;
use work.test_top_pkg.all;

-- Entity
entity test_top is
  port (
    -- AXI-Stream Bus for Ports
    s_axis_myinput_aclk     : in  std_logic;
    s_axis_myinput_aresetn  : in  std_logic;
    s_axis_myinput_tvalid   : in  std_logic;
    s_axis_myinput_tlast    : in  std_logic;
    s_axis_myinput_tdata    : in  std_logic_vector(PORTS_WIDTH-1 downto 0);
    m_axis_myoutput_aclk    : in  std_logic;
    m_axis_myoutput_aresetn : in  std_logic;
    m_axis_myoutput_tvalid  : out std_logic;
    m_axis_myoutput_tlast   : out std_logic;
    m_axis_myoutput_tdata   : out std_logic_vector(PORTS_WIDTH-1 downto 0);
    s_axis_test_in_aclk     : in  std_logic;
    s_axis_test_in_aresetn  : in  std_logic;
    s_axis_test_in_tready   : out std_logic;
    s_axis_test_in_tdata    : in  std_logic_vector(160-1 downto 0);
    s_axis_test_in_tuser    : in  std_logic_vector(128-1 downto 0);
    s_axis_test_in_tvalid   : in  std_logic;
    s_axis_test_in_tlast    : in  std_logic;
    m_axis_test_out_aclk    : in  std_logic;
    m_axis_test_out_aresetn : in  std_logic;
    m_axis_test_out_tready  : in  std_logic;
    m_axis_test_out_tdata   : out std_logic_vector(160-1 downto 0);
    m_axis_test_out_tuser   : out std_logic_vector(128-1 downto 0);
    m_axis_test_out_tvalid  : out std_logic;
    m_axis_test_out_tlast   : out std_logic;
    -- AXI4-Lite Bus for Properties
    S_AXI_ACLK             : in  std_logic;
    S_AXI_ARESETN          : in  std_logic;
    S_AXI_AWADDR           : in  std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
    S_AXI_AWPROT           : in  std_logic_vector(2 downto 0);
    S_AXI_AWVALID          : in  std_logic;
    S_AXI_AWREADY          : out std_logic;
    S_AXI_WDATA            : in  std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
    S_AXI_WSTRB            : in  std_logic_vector((PROPS_DATA_WIDTH/8)-1 downto 0);
    S_AXI_WVALID           : in  std_logic;
    S_AXI_WREADY           : out std_logic;
    S_AXI_BRESP            : out std_logic_vector(1 downto 0);
    S_AXI_BVALID           : out std_logic;
    S_AXI_BREADY           : in  std_logic;
    S_AXI_ARADDR           : in  std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
    S_AXI_ARPROT           : in  std_logic_vector(2 downto 0);
    S_AXI_ARVALID          : in  std_logic;
    S_AXI_ARREADY          : out std_logic;
    S_AXI_RDATA            : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
    S_AXI_RRESP            : out std_logic_vector(1 downto 0);
    S_AXI_RVALID           : out std_logic;
    S_AXI_RREADY           : in  std_logic;
    S_AXI_MIDDLE_ACLK      : in  std_logic;
    S_AXI_MIDDLE_ARESETN   : in  std_logic;
    S_AXI_MIDDLE_AWADDR    : in  std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
    S_AXI_MIDDLE_AWPROT    : in  std_logic_vector(2 downto 0);
    S_AXI_MIDDLE_AWVALID   : in  std_logic;
    S_AXI_MIDDLE_AWREADY   : out std_logic;
    S_AXI_MIDDLE_WDATA     : in  std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
    S_AXI_MIDDLE_WSTRB     : in  std_logic_vector((PROPS_DATA_WIDTH/8)-1 downto 0);
    S_AXI_MIDDLE_WVALID    : in  std_logic;
    S_AXI_MIDDLE_WREADY    : out std_logic;
    S_AXI_MIDDLE_BRESP     : out std_logic_vector(1 downto 0);
    S_AXI_MIDDLE_BVALID    : out std_logic;
    S_AXI_MIDDLE_BREADY    : in  std_logic;
    S_AXI_MIDDLE_ARADDR    : in  std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
    S_AXI_MIDDLE_ARPROT    : in  std_logic_vector(2 downto 0);
    S_AXI_MIDDLE_ARVALID   : in  std_logic;
    S_AXI_MIDDLE_ARREADY   : out std_logic;
    S_AXI_MIDDLE_RDATA     : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
    S_AXI_MIDDLE_RRESP     : out std_logic_vector(1 downto 0);
    S_AXI_MIDDLE_RVALID    : out std_logic;
    S_AXI_MIDDLE_RREADY    : in  std_logic;
    -- Sub-ip Software Configuration Bus
    s_swconfig_clk         : in  std_logic;
    s_swconfig_reset       : in  std_logic;
    s_swconfig_address     : in  std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
    s_swconfig_wr_enable   : in  std_logic;
    s_swconfig_wr_data     : in  std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
    s_swconfig_rd_enable   : in  std_logic;
    s_swconfig_rd_valid    : out std_logic;
    s_swconfig_rd_data     : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0)
  );
end entity test_top;

-- Architecture
architecture mixed of test_top is

  --------------------------------------------------------------------------------
  -- Constants
  --------------------------------------------------------------------------------
  constant TEST_RAM_ADDR_WIDTH : natural := integer(ceil(log2(real(TEST_RAM_DEPTH))));

  --------------------------------------------------------------------------------
  -- Components
  --------------------------------------------------------------------------------
  -- Autogenerated FINS HDL
  component test_top_axilite is
    generic (
      G_AXI_BYTE_INDEXED : boolean := True;
      G_AXI_ADDR_WIDTH   : natural := PROPS_ADDR_WIDTH;
      G_AXI_DATA_WIDTH   : natural := PROPS_DATA_WIDTH
    );
    port (
      -- AXI4-Lite Bus
      S_AXI_ACLK     : in  std_logic;
      S_AXI_ARESETN  : in  std_logic;
      S_AXI_AWADDR   : in  std_logic_vector(G_AXI_ADDR_WIDTH-1 downto 0);
      S_AXI_AWPROT   : in  std_logic_vector(2 downto 0);
      S_AXI_AWVALID  : in  std_logic;
      S_AXI_AWREADY  : out std_logic;
      S_AXI_WDATA    : in  std_logic_vector(G_AXI_DATA_WIDTH-1 downto 0);
      S_AXI_WSTRB    : in  std_logic_vector((G_AXI_DATA_WIDTH/8)-1 downto 0);
      S_AXI_WVALID   : in  std_logic;
      S_AXI_WREADY   : out std_logic;
      S_AXI_BRESP    : out std_logic_vector(1 downto 0);
      S_AXI_BVALID   : out std_logic;
      S_AXI_BREADY   : in  std_logic;
      S_AXI_ARADDR   : in  std_logic_vector(G_AXI_ADDR_WIDTH-1 downto 0);
      S_AXI_ARPROT   : in  std_logic_vector(2 downto 0);
      S_AXI_ARVALID  : in  std_logic;
      S_AXI_ARREADY  : out std_logic;
      S_AXI_RDATA    : out std_logic_vector(G_AXI_DATA_WIDTH-1 downto 0);
      S_AXI_RRESP    : out std_logic_vector(1 downto 0);
      S_AXI_RVALID   : out std_logic;
      S_AXI_RREADY   : in  std_logic;
      props_control  : out t_test_top_props_control;
      props_status   : in  t_test_top_props_status
    );
  end component;

  -- Autogenerated FINS HDL
  component test_top_axis is
    port (
      -- Input Port: myinput
      s_axis_myinput_aclk    : in  std_logic;
      s_axis_myinput_aresetn : in  std_logic;
      s_axis_myinput_tdata   : in  std_logic_vector(PORTS_WIDTH-1 downto 0);
      s_axis_myinput_tvalid  : in  std_logic;
      s_axis_myinput_tlast   : in  std_logic;
      -- Output Port: myoutput
      m_axis_myoutput_aclk    : in  std_logic;
      m_axis_myoutput_aresetn : in  std_logic;
      m_axis_myoutput_tdata   : out std_logic_vector(PORTS_WIDTH-1 downto 0);
      m_axis_myoutput_tvalid  : out std_logic;
      m_axis_myoutput_tlast   : out std_logic;
      -- Input Port: test_in
      s_axis_test_in_aclk    : in  std_logic;
      s_axis_test_in_aresetn : in  std_logic;
      s_axis_test_in_tready  : out std_logic;
      s_axis_test_in_tdata   : in  std_logic_vector(160-1 downto 0);
      s_axis_test_in_tuser   : in  std_logic_vector(128-1 downto 0);
      s_axis_test_in_tvalid  : in  std_logic;
      s_axis_test_in_tlast   : in  std_logic;
      -- Output Port: test_out
      m_axis_test_out_aclk    : in  std_logic;
      m_axis_test_out_aresetn : in  std_logic;
      m_axis_test_out_tready  : in  std_logic;
      m_axis_test_out_tdata   : out std_logic_vector(160-1 downto 0);
      m_axis_test_out_tuser   : out std_logic_vector(128-1 downto 0);
      m_axis_test_out_tvalid  : out std_logic;
      m_axis_test_out_tlast   : out std_logic;
      ports_in  : out t_test_top_ports_in;
      ports_out : in  t_test_top_ports_out
    );
  end component;

  -- Xilinx IP created by external_property_fifo.tcl script
  component xilinx_external_property_fifo
    port (
      clk   : in  std_logic;
      srst  : in  std_logic;
      din   : in  std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      wr_en : in  std_logic;
      rd_en : in  std_logic;
      dout  : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      full  : out std_logic;
      empty : out std_logic
    );
  end component;

  -- Xilinx IP created by memmap_property_ram.tcl script
  component xilinx_memmap_property_ram
    port (
      clka  : in std_logic;
      ena   : in std_logic;
      wea   : in std_logic_vector(0 downto 0);
      addra : in std_logic_vector(TEST_RAM_ADDR_WIDTH-1 downto 0);
      dina  : in std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      clkb  : in std_logic;
      enb   : in std_logic;
      addrb : in std_logic_vector(TEST_RAM_ADDR_WIDTH-1 downto 0);
      doutb : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0)
    );
  end component;

  -- Intel IP created by external_property_fifo.tcl script
  component intel_external_property_fifo is
    port (
      data  : in  std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      wrreq : in  std_logic;
      rdreq : in  std_logic;
      clock : in  std_logic;
      q     : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      full  : out std_logic;
      empty : out std_logic
    );
  end component;

  -- Intel IP created by memmap_property_ram.tcl script
  component intel_memmap_property_ram is
    port (
      data      : in  std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      q         : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      wraddress : in  std_logic_vector(TEST_RAM_ADDR_WIDTH-1 downto 0);
      rdaddress : in  std_logic_vector(TEST_RAM_ADDR_WIDTH-1 downto 0);
      wren      : in  std_logic;
      clock     : in  std_logic
    );
  end component;

  -- Sub-ip
  component test_middle_0 is
    port (
      -- AXI-Stream Bus for Ports
      s_axis_myinput_aclk     : in  std_logic;
      s_axis_myinput_aresetn  : in  std_logic;
      s_axis_myinput_tvalid   : in  std_logic;
      s_axis_myinput_tlast    : in  std_logic;
      s_axis_myinput_tdata    : in  std_logic_vector(PORTS_WIDTH-1 downto 0);
      m_axis_myoutput_aclk    : in  std_logic;
      m_axis_myoutput_aresetn : in  std_logic;
      m_axis_myoutput_tvalid  : out std_logic;
      m_axis_myoutput_tlast   : out std_logic;
      m_axis_myoutput_tdata   : out std_logic_vector(PORTS_WIDTH-1 downto 0);
      s_axis_test_in_aclk     : in  std_logic;
      s_axis_test_in_aresetn  : in  std_logic;
      s_axis_test_in_tready   : out std_logic;
      s_axis_test_in_tdata    : in  std_logic_vector(160-1 downto 0);
      s_axis_test_in_tuser    : in  std_logic_vector(128-1 downto 0);
      s_axis_test_in_tvalid   : in  std_logic;
      s_axis_test_in_tlast    : in  std_logic;
      m_axis_test_out_aclk    : in  std_logic;
      m_axis_test_out_aresetn : in  std_logic;
      m_axis_test_out_tready  : in  std_logic;
      m_axis_test_out_tdata   : out std_logic_vector(160-1 downto 0);
      m_axis_test_out_tuser   : out std_logic_vector(128-1 downto 0);
      m_axis_test_out_tvalid  : out std_logic;
      m_axis_test_out_tlast   : out std_logic;
      -- AXI4-Lite Bus for Properties
      S_AXI_ACLK             : in  std_logic;
      S_AXI_ARESETN          : in  std_logic;
      S_AXI_AWADDR           : in  std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
      S_AXI_AWPROT           : in  std_logic_vector(2 downto 0);
      S_AXI_AWVALID          : in  std_logic;
      S_AXI_AWREADY          : out std_logic;
      S_AXI_WDATA            : in  std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      S_AXI_WSTRB            : in  std_logic_vector((PROPS_DATA_WIDTH/8)-1 downto 0);
      S_AXI_WVALID           : in  std_logic;
      S_AXI_WREADY           : out std_logic;
      S_AXI_BRESP            : out std_logic_vector(1 downto 0);
      S_AXI_BVALID           : out std_logic;
      S_AXI_BREADY           : in  std_logic;
      S_AXI_ARADDR           : in  std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
      S_AXI_ARPROT           : in  std_logic_vector(2 downto 0);
      S_AXI_ARVALID          : in  std_logic;
      S_AXI_ARREADY          : out std_logic;
      S_AXI_RDATA            : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      S_AXI_RRESP            : out std_logic_vector(1 downto 0);
      S_AXI_RVALID           : out std_logic;
      S_AXI_RREADY           : in  std_logic;
      -- Sub-ip Software Configuration Bus
      s_swconfig_clk         : in  std_logic;
      s_swconfig_reset       : in  std_logic;
      s_swconfig_address     : in  std_logic_vector(PROPS_ADDR_WIDTH-1 downto 0);
      s_swconfig_wr_enable   : in  std_logic;
      s_swconfig_wr_data     : in  std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
      s_swconfig_rd_enable   : in  std_logic;
      s_swconfig_rd_valid    : out std_logic;
      s_swconfig_rd_data     : out std_logic_vector(PROPS_DATA_WIDTH-1 downto 0)
    );
  end component;

  --------------------------------------------------------------------------------
  -- Signals
  --------------------------------------------------------------------------------
  signal S_AXI_ARESET                 : std_logic;
  signal props_control                : t_test_top_props_control;
  signal props_status                 : t_test_top_props_status;
  signal external_property_register   : std_logic_vector(props_control.test_prop_write_only_external.wr_data'length-1 downto 0);
  signal memmap_property_ram_wr_en    : std_logic_vector(0 downto 0);
  signal memmap_property_ram_rd_en_q  : std_logic;
  signal memmap_property_ram_rd_en_qq : std_logic;
  signal memmap_property_register     : std_logic_vector(PROPS_DATA_WIDTH-1 downto 0);
  signal external_property_fifo_rd_en : std_logic;
  signal myinput_valid                : std_logic;
  signal myinput_last                 : std_logic;
  signal myinput_data                 : unsigned(PORTS_WIDTH-1 downto 0);
  signal myinput_valid_q              : std_logic;
  signal myinput_last_q               : std_logic;
  signal myinput_data_q               : unsigned(PORTS_WIDTH-1 downto 0);
  signal myoutput_valid               : std_logic;
  signal myoutput_last                : std_logic;
  signal myoutput_data                : std_logic_vector(PORTS_WIDTH-1 downto 0);
  signal test_out_tready              : std_logic;
  signal test_out_tdata               : std_logic_vector(160-1 downto 0);
  signal test_out_tuser               : std_logic_vector(128-1 downto 0);
  signal test_out_tvalid              : std_logic;
  signal test_out_tlast               : std_logic;
  signal ports_in                     : t_test_top_ports_in;
  signal ports_out                    : t_test_top_ports_out;

begin

  -- Invert reset for FIFO
  S_AXI_ARESET <= not S_AXI_ARESETN;

  --------------------------------------------------------------------------------
  -- Ports
  --------------------------------------------------------------------------------
  -- Instantiate ports module
  u_ports : test_top_axis
    port map (
      s_axis_myinput_aclk     => s_axis_myinput_aclk     ,
      s_axis_myinput_aresetn  => s_axis_myinput_aresetn  ,
      s_axis_myinput_tdata    => s_axis_myinput_tdata    ,
      s_axis_myinput_tvalid   => s_axis_myinput_tvalid   ,
      s_axis_myinput_tlast    => s_axis_myinput_tlast    ,
      m_axis_myoutput_aclk    => m_axis_myoutput_aclk    ,
      m_axis_myoutput_aresetn => m_axis_myoutput_aresetn ,
      m_axis_myoutput_tdata   => m_axis_myoutput_tdata   ,
      m_axis_myoutput_tvalid  => m_axis_myoutput_tvalid  ,
      m_axis_myoutput_tlast   => m_axis_myoutput_tlast   ,
      s_axis_test_in_aclk     => s_axis_test_in_aclk     ,
      s_axis_test_in_aresetn  => s_axis_test_in_aresetn  ,
      s_axis_test_in_tready   => s_axis_test_in_tready   ,
      s_axis_test_in_tdata    => s_axis_test_in_tdata    ,
      s_axis_test_in_tuser    => s_axis_test_in_tuser    ,
      s_axis_test_in_tvalid   => s_axis_test_in_tvalid   ,
      s_axis_test_in_tlast    => s_axis_test_in_tlast    ,
      m_axis_test_out_aclk    => m_axis_test_out_aclk    ,
      m_axis_test_out_aresetn => m_axis_test_out_aresetn ,
      m_axis_test_out_tready  => m_axis_test_out_tready  ,
      m_axis_test_out_tdata   => m_axis_test_out_tdata   ,
      m_axis_test_out_tuser   => m_axis_test_out_tuser   ,
      m_axis_test_out_tvalid  => m_axis_test_out_tvalid  ,
      m_axis_test_out_tlast   => m_axis_test_out_tlast   ,
      ports_in                => ports_in                ,
      ports_out               => ports_out               
    );

  --------------------------------------------------------------------------------
  -- Data Processing
  --------------------------------------------------------------------------------
  -- Synchronous process for data processsing
  s_data_processing : process (s_axis_myinput_aclk)
  begin
    if (rising_edge(s_axis_myinput_aclk)) then
      -- Data pipelines
      myinput_data <= ports_in.myinput.data;
      myinput_data_q <= resize(
        unsigned(myinput_data) * to_unsigned(TEST_PARAM_INTEGER, myinput_data'length),
        myinput_data'length
      );
      -- Control pipelines
      if (s_axis_myinput_aresetn = '0') then
        myinput_valid   <= '0';
        myinput_last    <= '0';
        myinput_valid_q <= '0';
        myinput_last_q  <= '0';
      else
        myinput_valid   <= ports_in.myinput.valid;
        myinput_last    <= ports_in.myinput.last;
        myinput_valid_q <= myinput_valid;
        myinput_last_q  <= myinput_last;
      end if;
    end if;
  end process s_data_processing;

  -- Instantiate sub-ip
  u_test_middle : test_middle_0
    port map (
      s_axis_myinput_aclk     => s_axis_myinput_aclk,
      s_axis_myinput_aresetn  => s_axis_myinput_aresetn,
      s_axis_myinput_tvalid   => myinput_valid_q,
      s_axis_myinput_tlast    => myinput_last_q,
      s_axis_myinput_tdata    => std_logic_vector(myinput_data_q),
      m_axis_myoutput_aclk    => m_axis_myoutput_aclk,
      m_axis_myoutput_aresetn => m_axis_myoutput_aresetn,
      m_axis_myoutput_tvalid  => myoutput_valid,
      m_axis_myoutput_tlast   => myoutput_last,
      m_axis_myoutput_tdata   => myoutput_data,
      s_axis_test_in_aclk     => s_axis_test_in_aclk,
      s_axis_test_in_aresetn  => s_axis_test_in_aresetn,
      s_axis_test_in_tready   => ports_out.test_in.ready,
      s_axis_test_in_tdata    => f_serialize_test_top_test_in_data(ports_in.test_in.data),
      s_axis_test_in_tuser    => f_serialize_test_top_test_in_metadata(ports_in.test_in.metadata),
      s_axis_test_in_tvalid   => ports_in.test_in.valid,
      s_axis_test_in_tlast    => ports_in.test_in.last,
      m_axis_test_out_aclk    => m_axis_test_out_aclk,
      m_axis_test_out_aresetn => m_axis_test_out_aresetn,
      m_axis_test_out_tready  => test_out_tready,
      m_axis_test_out_tdata   => test_out_tdata,
      m_axis_test_out_tuser   => test_out_tuser,
      m_axis_test_out_tvalid  => test_out_tvalid,
      m_axis_test_out_tlast   => test_out_tlast,
      S_AXI_ACLK              => S_AXI_MIDDLE_ACLK,
      S_AXI_ARESETN           => S_AXI_MIDDLE_ARESETN,
      S_AXI_AWADDR            => S_AXI_MIDDLE_AWADDR,
      S_AXI_AWPROT            => S_AXI_MIDDLE_AWPROT,
      S_AXI_AWVALID           => S_AXI_MIDDLE_AWVALID,
      S_AXI_AWREADY           => S_AXI_MIDDLE_AWREADY,
      S_AXI_WDATA             => S_AXI_MIDDLE_WDATA,
      S_AXI_WSTRB             => S_AXI_MIDDLE_WSTRB,
      S_AXI_WVALID            => S_AXI_MIDDLE_WVALID,
      S_AXI_WREADY            => S_AXI_MIDDLE_WREADY,
      S_AXI_BRESP             => S_AXI_MIDDLE_BRESP,
      S_AXI_BVALID            => S_AXI_MIDDLE_BVALID,
      S_AXI_BREADY            => S_AXI_MIDDLE_BREADY,
      S_AXI_ARADDR            => S_AXI_MIDDLE_ARADDR,
      S_AXI_ARPROT            => S_AXI_MIDDLE_ARPROT,
      S_AXI_ARVALID           => S_AXI_MIDDLE_ARVALID,
      S_AXI_ARREADY           => S_AXI_MIDDLE_ARREADY,
      S_AXI_RDATA             => S_AXI_MIDDLE_RDATA,
      S_AXI_RRESP             => S_AXI_MIDDLE_RRESP,
      S_AXI_RVALID            => S_AXI_MIDDLE_RVALID,
      S_AXI_RREADY            => S_AXI_MIDDLE_RREADY,
      s_swconfig_clk          => s_swconfig_clk,
      s_swconfig_reset        => s_swconfig_reset,
      s_swconfig_address      => s_swconfig_address,
      s_swconfig_wr_enable    => s_swconfig_wr_enable,
      s_swconfig_wr_data      => s_swconfig_wr_data,
      s_swconfig_rd_enable    => s_swconfig_rd_enable,
      s_swconfig_rd_valid     => s_swconfig_rd_valid,
      s_swconfig_rd_data      => s_swconfig_rd_data
    );

  -- Assign output ports
  ports_out.myoutput.valid    <= myoutput_valid;
  ports_out.myoutput.last     <= myoutput_last;
  ports_out.myoutput.data     <= f_unserialize_test_top_myoutput_data(myoutput_data);
  ports_out.test_out.data     <= f_unserialize_test_top_test_out_data(test_out_tdata);
  ports_out.test_out.metadata <= f_unserialize_test_top_test_out_metadata(test_out_tuser);
  ports_out.test_out.valid    <= test_out_tvalid;
  ports_out.test_out.last     <= test_out_tlast;
  test_out_tready             <= ports_in.test_out.ready;

  --------------------------------------------------------------------------------
  -- Properties
  --------------------------------------------------------------------------------
  -- Instantiate the auto-generated AXI4-Lite module
  u_properties : test_top_axilite
    port map (
      S_AXI_ACLK    => S_AXI_ACLK    ,
      S_AXI_ARESETN => S_AXI_ARESETN ,
      S_AXI_AWADDR  => S_AXI_AWADDR  ,
      S_AXI_AWPROT  => S_AXI_AWPROT  ,
      S_AXI_AWVALID => S_AXI_AWVALID ,
      S_AXI_AWREADY => S_AXI_AWREADY ,
      S_AXI_WDATA   => S_AXI_WDATA   ,
      S_AXI_WSTRB   => S_AXI_WSTRB   ,
      S_AXI_WVALID  => S_AXI_WVALID  ,
      S_AXI_WREADY  => S_AXI_WREADY  ,
      S_AXI_BRESP   => S_AXI_BRESP   ,
      S_AXI_BVALID  => S_AXI_BVALID  ,
      S_AXI_BREADY  => S_AXI_BREADY  ,
      S_AXI_ARADDR  => S_AXI_ARADDR  ,
      S_AXI_ARPROT  => S_AXI_ARPROT  ,
      S_AXI_ARVALID => S_AXI_ARVALID ,
      S_AXI_ARREADY => S_AXI_ARREADY ,
      S_AXI_RDATA   => S_AXI_RDATA   ,
      S_AXI_RRESP   => S_AXI_RRESP   ,
      S_AXI_RVALID  => S_AXI_RVALID  ,
      S_AXI_RREADY  => S_AXI_RREADY  ,
      props_control => props_control ,
      props_status  => props_status  
    );

  --------------------------------------------------------------------------------
  -- Testing elements for "read-write-external"
  --------------------------------------------------------------------------------
  -- FWFT FIFO instantitation for test
  u_gen_xilinx_external_property_fifo : if (USE_XILINX) generate
    u_external_property_fifo : xilinx_external_property_fifo
      port map (
        clk   => s_swconfig_clk,
        srst  => s_swconfig_reset,
        din   => props_control.test_prop_read_write_external.wr_data,
        wr_en => props_control.test_prop_read_write_external.wr_en,
        rd_en => external_property_fifo_rd_en,
        dout  => props_status.test_prop_read_write_external.rd_data,
        full  => open,
        empty => open
      );
  end generate u_gen_xilinx_external_property_fifo;
  u_gen_intel_external_property_fifo : if (not USE_XILINX) generate
    u_external_property_fifo : intel_external_property_fifo
      port map (
        clock   => s_swconfig_clk,
        data    => props_control.test_prop_read_write_external.wr_data,
        wrreq   => props_control.test_prop_read_write_external.wr_en,
        rdreq   => external_property_fifo_rd_en,
        q       => props_status.test_prop_read_write_external.rd_data,
        full    => open,
        empty   => open
      );
  end generate u_gen_intel_external_property_fifo;

  -- Synchronous process to delay the fifo read enable one clock just due to this FIFO's timing
  s_external_property_fifo : process(s_swconfig_clk)
  begin
    if (rising_edge(s_swconfig_clk)) then
      if (s_swconfig_reset = '1') then
        external_property_fifo_rd_en <= '0';
      else
        external_property_fifo_rd_en <= props_control.test_prop_read_write_external.rd_en;
      end if;
    end if;
  end process s_external_property_fifo;

  -- Since this is a FWFT FIFO, the read data is valid as soon as the FIFO is read
  props_status.test_prop_read_write_external.rd_valid <= props_control.test_prop_read_write_external.rd_en;

  --------------------------------------------------------------------------------
  -- Testing elements for "write-only-external" and "read-only-external"
  --------------------------------------------------------------------------------
  -- Synchronous process for external property write
  s_external_property_register : process(S_AXI_ACLK)
  begin
    if (rising_edge(S_AXI_ACLK)) then
      if (S_AXI_ARESETN = '0') then
        external_property_register <= (others => '0');
      else
        if (props_control.test_prop_write_only_external.wr_en = '1') then
          external_property_register <= props_control.test_prop_write_only_external.wr_data;
        end if;
      end if;
    end if;
  end process s_external_property_register;

  -- Assign read signals to register written above
  props_status.test_prop_read_only_external.rd_valid <= props_control.test_prop_read_only_external.rd_en;
  props_status.test_prop_read_only_external.rd_data  <= external_property_register;

  --------------------------------------------------------------------------------
  -- Testing elements for "read-write-memmap"
  --------------------------------------------------------------------------------
  -- Simple Dual Port RAM for test
  u_gen_xilinx_memmap_property_ram : if (USE_XILINX) generate
    u_memmap_property_ram : xilinx_memmap_property_ram
      port map (
        clka  => s_swconfig_clk,
        ena   => '1',
        wea   => memmap_property_ram_wr_en,
        addra => props_control.test_prop_read_write_memmap.wr_addr,
        dina  => props_control.test_prop_read_write_memmap.wr_data,
        clkb  => s_swconfig_clk,
        enb   => '1',
        addrb => props_control.test_prop_read_write_memmap.rd_addr,
        doutb => props_status.test_prop_read_write_memmap.rd_data
      );
  end generate u_gen_xilinx_memmap_property_ram;
  u_gen_intel_memmap_property_ram : if (not USE_XILINX) generate
    u_memmap_property_ram : intel_memmap_property_ram
      port map (
        clock     => s_swconfig_clk,
        wren      => props_control.test_prop_read_write_memmap.wr_en,
        wraddress => props_control.test_prop_read_write_memmap.wr_addr,
        data      => props_control.test_prop_read_write_memmap.wr_data,
        rdaddress => props_control.test_prop_read_write_memmap.rd_addr,
        q         => props_status.test_prop_read_write_memmap.rd_data
      );
  end generate u_gen_intel_memmap_property_ram;

  -- Remap the write enable to a std_logic_vector of width 1
  memmap_property_ram_wr_en(0) <= props_control.test_prop_read_write_memmap.wr_en;

  -- Synchronous process to delay the read enable 2 clocks
  s_memmap_property_ram : process (S_AXI_ACLK)
  begin
    if (rising_edge(S_AXI_ACLK)) then
      if (S_AXI_ARESETN = '0') then
        memmap_property_ram_rd_en_q  <= '0';
        memmap_property_ram_rd_en_qq <= '0';
      else
        memmap_property_ram_rd_en_q  <= props_control.test_prop_read_write_memmap.rd_en;
        memmap_property_ram_rd_en_qq <= memmap_property_ram_rd_en_q;
      end if;
    end if;
  end process s_memmap_property_ram;

  -- Assign the read valid to the delayed copy of the read enable due to the latency of the
  -- Simple Dual Port RAM
  props_status.test_prop_read_write_memmap.rd_valid <= memmap_property_ram_rd_en_qq;

  --------------------------------------------------------------------------------
  -- Testing elements for "write-only-memmap" and "read-only-memmap"
  --------------------------------------------------------------------------------
  -- Note: Since this property has a length of 1, the addresses are unused and
  --       the behavior mirrors an "external" property. This use case is unusual
  --       but is tested for completeness.

  -- Synchronous process for memmap property write
  s_memmap_property_register : process(S_AXI_ACLK)
  begin
    if (rising_edge(S_AXI_ACLK)) then
      if (S_AXI_ARESETN = '0') then
        memmap_property_register <= (others => '0');
      else
        if (props_control.test_prop_write_only_memmap.wr_en = '1') then
          memmap_property_register <= props_control.test_prop_write_only_memmap.wr_data;
        end if;
      end if;
    end if;
  end process s_memmap_property_register;

  -- Assign read signals to register written above
  props_status.test_prop_read_only_memmap.rd_valid <= props_control.test_prop_read_only_memmap.rd_en;
  props_status.test_prop_read_only_memmap.rd_data  <= memmap_property_register;

  --------------------------------------------------------------------------------
  -- Testing elements for "read-only-data"
  --------------------------------------------------------------------------------
  props_status.test_prop_read_only_data(0).rd_data <= std_logic_vector(to_unsigned(0, PROPS_DATA_WIDTH));
  props_status.test_prop_read_only_data(1).rd_data <= std_logic_vector(to_unsigned(1, PROPS_DATA_WIDTH));
  props_status.test_prop_read_only_data(2).rd_data <= std_logic_vector(to_unsigned(2, PROPS_DATA_WIDTH));
  props_status.test_prop_read_only_data(3).rd_data <= std_logic_vector(to_unsigned(3, PROPS_DATA_WIDTH));

end mixed;
